
module pipelined_fir_filter (
    input wire clk,
    input wire rst,
    input wire signed [15:0] data_in,
    output reg signed [31:0] data_out
);

localparam TAPS = 100;
localparam signed [15:0] COEFF_0 = -16'sd5;
localparam signed [15:0] COEFF_1 = -16'sd14;
localparam signed [15:0] COEFF_2 = -16'sd18;
localparam signed [15:0] COEFF_3 = -16'sd16;
localparam signed [15:0] COEFF_4 = -16'sd6;
localparam signed [15:0] COEFF_5 = 16'sd7;
localparam signed [15:0] COEFF_6 = 16'sd21;
localparam signed [15:0] COEFF_7 = 16'sd30;
localparam signed [15:0] COEFF_8 = 16'sd28;
localparam signed [15:0] COEFF_9 = 16'sd12;
localparam signed [15:0] COEFF_10 = -16'sd13;
localparam signed [15:0] COEFF_11 = -16'sd41;
localparam signed [15:0] COEFF_12 = -16'sd57;
localparam signed [15:0] COEFF_13 = -16'sd52;
localparam signed [15:0] COEFF_14 = -16'sd22;
localparam signed [15:0] COEFF_15 = 16'sd25;
localparam signed [15:0] COEFF_16 = 16'sd75;
localparam signed [15:0] COEFF_17 = 16'sd103;
localparam signed [15:0] COEFF_18 = 16'sd93;
localparam signed [15:0] COEFF_19 = 16'sd39;
localparam signed [15:0] COEFF_20 = -16'sd44;
localparam signed [15:0] COEFF_21 = -16'sd127;
localparam signed [15:0] COEFF_22 = -16'sd174;
localparam signed [15:0] COEFF_23 = -16'sd155;
localparam signed [15:0] COEFF_24 = -16'sd65;
localparam signed [15:0] COEFF_25 = 16'sd72;
localparam signed [15:0] COEFF_26 = 16'sd207;
localparam signed [15:0] COEFF_27 = 16'sd281;
localparam signed [15:0] COEFF_28 = 16'sd249;
localparam signed [15:0] COEFF_29 = 16'sd104;
localparam signed [15:0] COEFF_30 = -16'sd114;
localparam signed [15:0] COEFF_31 = -16'sd327;
localparam signed [15:0] COEFF_32 = -16'sd444;
localparam signed [15:0] COEFF_33 = -16'sd394;
localparam signed [15:0] COEFF_34 = -16'sd165;
localparam signed [15:0] COEFF_35 = 16'sd182;
localparam signed [15:0] COEFF_36 = 16'sd526;
localparam signed [15:0] COEFF_37 = 16'sd720;
localparam signed [15:0] COEFF_38 = 16'sd648;
localparam signed [15:0] COEFF_39 = 16'sd277;
localparam signed [15:0] COEFF_40 = -16'sd312;
localparam signed [15:0] COEFF_41 = -16'sd929;
localparam signed [15:0] COEFF_42 = -16'sd1321;
localparam signed [15:0] COEFF_43 = -16'sd1250;
localparam signed [15:0] COEFF_44 = -16'sd570;
localparam signed [15:0] COEFF_45 = 16'sd704;
localparam signed [15:0] COEFF_46 = 16'sd2387;
localparam signed [15:0] COEFF_47 = 16'sd4154;
localparam signed [15:0] COEFF_48 = 16'sd5622;
localparam signed [15:0] COEFF_49 = 16'sd6454;
localparam signed [15:0] COEFF_50 = 16'sd6454;
localparam signed [15:0] COEFF_51 = 16'sd5622;
localparam signed [15:0] COEFF_52 = 16'sd4154;
localparam signed [15:0] COEFF_53 = 16'sd2387;
localparam signed [15:0] COEFF_54 = 16'sd704;
localparam signed [15:0] COEFF_55 = -16'sd570;
localparam signed [15:0] COEFF_56 = -16'sd1250;
localparam signed [15:0] COEFF_57 = -16'sd1321;
localparam signed [15:0] COEFF_58 = -16'sd929;
localparam signed [15:0] COEFF_59 = -16'sd312;
localparam signed [15:0] COEFF_60 = 16'sd277;
localparam signed [15:0] COEFF_61 = 16'sd648;
localparam signed [15:0] COEFF_62 = 16'sd720;
localparam signed [15:0] COEFF_63 = 16'sd526;
localparam signed [15:0] COEFF_64 = 16'sd182;
localparam signed [15:0] COEFF_65 = -16'sd165;
localparam signed [15:0] COEFF_66 = -16'sd394;
localparam signed [15:0] COEFF_67 = -16'sd444;
localparam signed [15:0] COEFF_68 = -16'sd327;
localparam signed [15:0] COEFF_69 = -16'sd114;
localparam signed [15:0] COEFF_70 = 16'sd104;
localparam signed [15:0] COEFF_71 = 16'sd249;
localparam signed [15:0] COEFF_72 = 16'sd281;
localparam signed [15:0] COEFF_73 = 16'sd207;
localparam signed [15:0] COEFF_74 = 16'sd72;
localparam signed [15:0] COEFF_75 = -16'sd65;
localparam signed [15:0] COEFF_76 = -16'sd155;
localparam signed [15:0] COEFF_77 = -16'sd174;
localparam signed [15:0] COEFF_78 = -16'sd127;
localparam signed [15:0] COEFF_79 = -16'sd44;
localparam signed [15:0] COEFF_80 = 16'sd39;
localparam signed [15:0] COEFF_81 = 16'sd93;
localparam signed [15:0] COEFF_82 = 16'sd103;
localparam signed [15:0] COEFF_83 = 16'sd75;
localparam signed [15:0] COEFF_84 = 16'sd25;
localparam signed [15:0] COEFF_85 = -16'sd22;
localparam signed [15:0] COEFF_86 = -16'sd52;
localparam signed [15:0] COEFF_87 = -16'sd57;
localparam signed [15:0] COEFF_88 = -16'sd41;
localparam signed [15:0] COEFF_89 = -16'sd13;
localparam signed [15:0] COEFF_90 = 16'sd12;
localparam signed [15:0] COEFF_91 = 16'sd28;
localparam signed [15:0] COEFF_92 = 16'sd30;
localparam signed [15:0] COEFF_93 = 16'sd21;
localparam signed [15:0] COEFF_94 = 16'sd7;
localparam signed [15:0] COEFF_95 = -16'sd6;
localparam signed [15:0] COEFF_96 = -16'sd16;
localparam signed [15:0] COEFF_97 = -16'sd18;
localparam signed [15:0] COEFF_98 = -16'sd14;
localparam signed [15:0] COEFF_99 = -16'sd5;

reg signed [15:0] shift_reg[TAPS-1:0];
reg signed [31:0] pipe_stage_0[0:0]; // Pipeline stage for COEFF_0
reg signed [31:0] pipe_stage_1[0:0]; // Pipeline stage for COEFF_1
reg signed [31:0] pipe_stage_2[0:0]; // Pipeline stage for COEFF_2
reg signed [31:0] pipe_stage_3[0:0]; // Pipeline stage for COEFF_3
reg signed [31:0] pipe_stage_4[0:0]; // Pipeline stage for COEFF_4
reg signed [31:0] pipe_stage_5[0:0]; // Pipeline stage for COEFF_5
reg signed [31:0] pipe_stage_6[0:0]; // Pipeline stage for COEFF_6
reg signed [31:0] pipe_stage_7[0:0]; // Pipeline stage for COEFF_7
reg signed [31:0] pipe_stage_8[0:0]; // Pipeline stage for COEFF_8
reg signed [31:0] pipe_stage_9[0:0]; // Pipeline stage for COEFF_9
reg signed [31:0] pipe_stage_10[0:0]; // Pipeline stage for COEFF_10
reg signed [31:0] pipe_stage_11[0:0]; // Pipeline stage for COEFF_11
reg signed [31:0] pipe_stage_12[0:0]; // Pipeline stage for COEFF_12
reg signed [31:0] pipe_stage_13[0:0]; // Pipeline stage for COEFF_13
reg signed [31:0] pipe_stage_14[0:0]; // Pipeline stage for COEFF_14
reg signed [31:0] pipe_stage_15[0:0]; // Pipeline stage for COEFF_15
reg signed [31:0] pipe_stage_16[0:0]; // Pipeline stage for COEFF_16
reg signed [31:0] pipe_stage_17[0:0]; // Pipeline stage for COEFF_17
reg signed [31:0] pipe_stage_18[0:0]; // Pipeline stage for COEFF_18
reg signed [31:0] pipe_stage_19[0:0]; // Pipeline stage for COEFF_19
reg signed [31:0] pipe_stage_20[0:0]; // Pipeline stage for COEFF_20
reg signed [31:0] pipe_stage_21[0:0]; // Pipeline stage for COEFF_21
reg signed [31:0] pipe_stage_22[0:0]; // Pipeline stage for COEFF_22
reg signed [31:0] pipe_stage_23[0:0]; // Pipeline stage for COEFF_23
reg signed [31:0] pipe_stage_24[0:0]; // Pipeline stage for COEFF_24
reg signed [31:0] pipe_stage_25[0:0]; // Pipeline stage for COEFF_25
reg signed [31:0] pipe_stage_26[0:0]; // Pipeline stage for COEFF_26
reg signed [31:0] pipe_stage_27[0:0]; // Pipeline stage for COEFF_27
reg signed [31:0] pipe_stage_28[0:0]; // Pipeline stage for COEFF_28
reg signed [31:0] pipe_stage_29[0:0]; // Pipeline stage for COEFF_29
reg signed [31:0] pipe_stage_30[0:0]; // Pipeline stage for COEFF_30
reg signed [31:0] pipe_stage_31[0:0]; // Pipeline stage for COEFF_31
reg signed [31:0] pipe_stage_32[0:0]; // Pipeline stage for COEFF_32
reg signed [31:0] pipe_stage_33[0:0]; // Pipeline stage for COEFF_33
reg signed [31:0] pipe_stage_34[0:0]; // Pipeline stage for COEFF_34
reg signed [31:0] pipe_stage_35[0:0]; // Pipeline stage for COEFF_35
reg signed [31:0] pipe_stage_36[0:0]; // Pipeline stage for COEFF_36
reg signed [31:0] pipe_stage_37[0:0]; // Pipeline stage for COEFF_37
reg signed [31:0] pipe_stage_38[0:0]; // Pipeline stage for COEFF_38
reg signed [31:0] pipe_stage_39[0:0]; // Pipeline stage for COEFF_39
reg signed [31:0] pipe_stage_40[0:0]; // Pipeline stage for COEFF_40
reg signed [31:0] pipe_stage_41[0:0]; // Pipeline stage for COEFF_41
reg signed [31:0] pipe_stage_42[0:0]; // Pipeline stage for COEFF_42
reg signed [31:0] pipe_stage_43[0:0]; // Pipeline stage for COEFF_43
reg signed [31:0] pipe_stage_44[0:0]; // Pipeline stage for COEFF_44
reg signed [31:0] pipe_stage_45[0:0]; // Pipeline stage for COEFF_45
reg signed [31:0] pipe_stage_46[0:0]; // Pipeline stage for COEFF_46
reg signed [31:0] pipe_stage_47[0:0]; // Pipeline stage for COEFF_47
reg signed [31:0] pipe_stage_48[0:0]; // Pipeline stage for COEFF_48
reg signed [31:0] pipe_stage_49[0:0]; // Pipeline stage for COEFF_49
reg signed [31:0] pipe_stage_50[0:0]; // Pipeline stage for COEFF_50
reg signed [31:0] pipe_stage_51[0:0]; // Pipeline stage for COEFF_51
reg signed [31:0] pipe_stage_52[0:0]; // Pipeline stage for COEFF_52
reg signed [31:0] pipe_stage_53[0:0]; // Pipeline stage for COEFF_53
reg signed [31:0] pipe_stage_54[0:0]; // Pipeline stage for COEFF_54
reg signed [31:0] pipe_stage_55[0:0]; // Pipeline stage for COEFF_55
reg signed [31:0] pipe_stage_56[0:0]; // Pipeline stage for COEFF_56
reg signed [31:0] pipe_stage_57[0:0]; // Pipeline stage for COEFF_57
reg signed [31:0] pipe_stage_58[0:0]; // Pipeline stage for COEFF_58
reg signed [31:0] pipe_stage_59[0:0]; // Pipeline stage for COEFF_59
reg signed [31:0] pipe_stage_60[0:0]; // Pipeline stage for COEFF_60
reg signed [31:0] pipe_stage_61[0:0]; // Pipeline stage for COEFF_61
reg signed [31:0] pipe_stage_62[0:0]; // Pipeline stage for COEFF_62
reg signed [31:0] pipe_stage_63[0:0]; // Pipeline stage for COEFF_63
reg signed [31:0] pipe_stage_64[0:0]; // Pipeline stage for COEFF_64
reg signed [31:0] pipe_stage_65[0:0]; // Pipeline stage for COEFF_65
reg signed [31:0] pipe_stage_66[0:0]; // Pipeline stage for COEFF_66
reg signed [31:0] pipe_stage_67[0:0]; // Pipeline stage for COEFF_67
reg signed [31:0] pipe_stage_68[0:0]; // Pipeline stage for COEFF_68
reg signed [31:0] pipe_stage_69[0:0]; // Pipeline stage for COEFF_69
reg signed [31:0] pipe_stage_70[0:0]; // Pipeline stage for COEFF_70
reg signed [31:0] pipe_stage_71[0:0]; // Pipeline stage for COEFF_71
reg signed [31:0] pipe_stage_72[0:0]; // Pipeline stage for COEFF_72
reg signed [31:0] pipe_stage_73[0:0]; // Pipeline stage for COEFF_73
reg signed [31:0] pipe_stage_74[0:0]; // Pipeline stage for COEFF_74
reg signed [31:0] pipe_stage_75[0:0]; // Pipeline stage for COEFF_75
reg signed [31:0] pipe_stage_76[0:0]; // Pipeline stage for COEFF_76
reg signed [31:0] pipe_stage_77[0:0]; // Pipeline stage for COEFF_77
reg signed [31:0] pipe_stage_78[0:0]; // Pipeline stage for COEFF_78
reg signed [31:0] pipe_stage_79[0:0]; // Pipeline stage for COEFF_79
reg signed [31:0] pipe_stage_80[0:0]; // Pipeline stage for COEFF_80
reg signed [31:0] pipe_stage_81[0:0]; // Pipeline stage for COEFF_81
reg signed [31:0] pipe_stage_82[0:0]; // Pipeline stage for COEFF_82
reg signed [31:0] pipe_stage_83[0:0]; // Pipeline stage for COEFF_83
reg signed [31:0] pipe_stage_84[0:0]; // Pipeline stage for COEFF_84
reg signed [31:0] pipe_stage_85[0:0]; // Pipeline stage for COEFF_85
reg signed [31:0] pipe_stage_86[0:0]; // Pipeline stage for COEFF_86
reg signed [31:0] pipe_stage_87[0:0]; // Pipeline stage for COEFF_87
reg signed [31:0] pipe_stage_88[0:0]; // Pipeline stage for COEFF_88
reg signed [31:0] pipe_stage_89[0:0]; // Pipeline stage for COEFF_89
reg signed [31:0] pipe_stage_90[0:0]; // Pipeline stage for COEFF_90
reg signed [31:0] pipe_stage_91[0:0]; // Pipeline stage for COEFF_91
reg signed [31:0] pipe_stage_92[0:0]; // Pipeline stage for COEFF_92
reg signed [31:0] pipe_stage_93[0:0]; // Pipeline stage for COEFF_93
reg signed [31:0] pipe_stage_94[0:0]; // Pipeline stage for COEFF_94
reg signed [31:0] pipe_stage_95[0:0]; // Pipeline stage for COEFF_95
reg signed [31:0] pipe_stage_96[0:0]; // Pipeline stage for COEFF_96
reg signed [31:0] pipe_stage_97[0:0]; // Pipeline stage for COEFF_97
reg signed [31:0] pipe_stage_98[0:0]; // Pipeline stage for COEFF_98
reg signed [31:0] pipe_stage_99[0:0]; // Pipeline stage for COEFF_99

integer i;

always @(posedge clk) begin
    if (rst) begin
        // Reset logic
        for (i = 0; i < TAPS; i = i + 1) begin
            shift_reg[i] <= 0;
        end
        data_out <= 0;
    end else begin
        // Shift the input data through the register
        for (i = TAPS-1; i > 0; i = i - 1) begin
            shift_reg[i] <= shift_reg[i - 1];
        end
        shift_reg[0] <= data_in;

        // Pipeline processing
        pipe_stage_0[0] = shift_reg[0] * COEFF_0;
        pipe_stage_1[0] = shift_reg[1] * COEFF_1;
        pipe_stage_2[0] = shift_reg[2] * COEFF_2;
        pipe_stage_3[0] = shift_reg[3] * COEFF_3;
        pipe_stage_4[0] = shift_reg[4] * COEFF_4;
        pipe_stage_5[0] = shift_reg[5] * COEFF_5;
        pipe_stage_6[0] = shift_reg[6] * COEFF_6;
        pipe_stage_7[0] = shift_reg[7] * COEFF_7;
        pipe_stage_8[0] = shift_reg[8] * COEFF_8;
        pipe_stage_9[0] = shift_reg[9] * COEFF_9;
        pipe_stage_10[0] = shift_reg[10] * COEFF_10;
        pipe_stage_11[0] = shift_reg[11] * COEFF_11;
        pipe_stage_12[0] = shift_reg[12] * COEFF_12;
        pipe_stage_13[0] = shift_reg[13] * COEFF_13;
        pipe_stage_14[0] = shift_reg[14] * COEFF_14;
        pipe_stage_15[0] = shift_reg[15] * COEFF_15;
        pipe_stage_16[0] = shift_reg[16] * COEFF_16;
        pipe_stage_17[0] = shift_reg[17] * COEFF_17;
        pipe_stage_18[0] = shift_reg[18] * COEFF_18;
        pipe_stage_19[0] = shift_reg[19] * COEFF_19;
        pipe_stage_20[0] = shift_reg[20] * COEFF_20;
        pipe_stage_21[0] = shift_reg[21] * COEFF_21;
        pipe_stage_22[0] = shift_reg[22] * COEFF_22;
        pipe_stage_23[0] = shift_reg[23] * COEFF_23;
        pipe_stage_24[0] = shift_reg[24] * COEFF_24;
        pipe_stage_25[0] = shift_reg[25] * COEFF_25;
        pipe_stage_26[0] = shift_reg[26] * COEFF_26;
        pipe_stage_27[0] = shift_reg[27] * COEFF_27;
        pipe_stage_28[0] = shift_reg[28] * COEFF_28;
        pipe_stage_29[0] = shift_reg[29] * COEFF_29;
        pipe_stage_30[0] = shift_reg[30] * COEFF_30;
        pipe_stage_31[0] = shift_reg[31] * COEFF_31;
        pipe_stage_32[0] = shift_reg[32] * COEFF_32;
        pipe_stage_33[0] = shift_reg[33] * COEFF_33;
        pipe_stage_34[0] = shift_reg[34] * COEFF_34;
        pipe_stage_35[0] = shift_reg[35] * COEFF_35;
        pipe_stage_36[0] = shift_reg[36] * COEFF_36;
        pipe_stage_37[0] = shift_reg[37] * COEFF_37;
        pipe_stage_38[0] = shift_reg[38] * COEFF_38;
        pipe_stage_39[0] = shift_reg[39] * COEFF_39;
        pipe_stage_40[0] = shift_reg[40] * COEFF_40;
        pipe_stage_41[0] = shift_reg[41] * COEFF_41;
        pipe_stage_42[0] = shift_reg[42] * COEFF_42;
        pipe_stage_43[0] = shift_reg[43] * COEFF_43;
        pipe_stage_44[0] = shift_reg[44] * COEFF_44;
        pipe_stage_45[0] = shift_reg[45] * COEFF_45;
        pipe_stage_46[0] = shift_reg[46] * COEFF_46;
        pipe_stage_47[0] = shift_reg[47] * COEFF_47;
        pipe_stage_48[0] = shift_reg[48] * COEFF_48;
        pipe_stage_49[0] = shift_reg[49] * COEFF_49;
        pipe_stage_50[0] = shift_reg[50] * COEFF_50;
        pipe_stage_51[0] = shift_reg[51] * COEFF_51;
        pipe_stage_52[0] = shift_reg[52] * COEFF_52;
        pipe_stage_53[0] = shift_reg[53] * COEFF_53;
        pipe_stage_54[0] = shift_reg[54] * COEFF_54;
        pipe_stage_55[0] = shift_reg[55] * COEFF_55;
        pipe_stage_56[0] = shift_reg[56] * COEFF_56;
        pipe_stage_57[0] = shift_reg[57] * COEFF_57;
        pipe_stage_58[0] = shift_reg[58] * COEFF_58;
        pipe_stage_59[0] = shift_reg[59] * COEFF_59;
        pipe_stage_60[0] = shift_reg[60] * COEFF_60;
        pipe_stage_61[0] = shift_reg[61] * COEFF_61;
        pipe_stage_62[0] = shift_reg[62] * COEFF_62;
        pipe_stage_63[0] = shift_reg[63] * COEFF_63;
        pipe_stage_64[0] = shift_reg[64] * COEFF_64;
        pipe_stage_65[0] = shift_reg[65] * COEFF_65;
        pipe_stage_66[0] = shift_reg[66] * COEFF_66;
        pipe_stage_67[0] = shift_reg[67] * COEFF_67;
        pipe_stage_68[0] = shift_reg[68] * COEFF_68;
        pipe_stage_69[0] = shift_reg[69] * COEFF_69;
        pipe_stage_70[0] = shift_reg[70] * COEFF_70;
        pipe_stage_71[0] = shift_reg[71] * COEFF_71;
        pipe_stage_72[0] = shift_reg[72] * COEFF_72;
        pipe_stage_73[0] = shift_reg[73] * COEFF_73;
        pipe_stage_74[0] = shift_reg[74] * COEFF_74;
        pipe_stage_75[0] = shift_reg[75] * COEFF_75;
        pipe_stage_76[0] = shift_reg[76] * COEFF_76;
        pipe_stage_77[0] = shift_reg[77] * COEFF_77;
        pipe_stage_78[0] = shift_reg[78] * COEFF_78;
        pipe_stage_79[0] = shift_reg[79] * COEFF_79;
        pipe_stage_80[0] = shift_reg[80] * COEFF_80;
        pipe_stage_81[0] = shift_reg[81] * COEFF_81;
        pipe_stage_82[0] = shift_reg[82] * COEFF_82;
        pipe_stage_83[0] = shift_reg[83] * COEFF_83;
        pipe_stage_84[0] = shift_reg[84] * COEFF_84;
        pipe_stage_85[0] = shift_reg[85] * COEFF_85;
        pipe_stage_86[0] = shift_reg[86] * COEFF_86;
        pipe_stage_87[0] = shift_reg[87] * COEFF_87;
        pipe_stage_88[0] = shift_reg[88] * COEFF_88;
        pipe_stage_89[0] = shift_reg[89] * COEFF_89;
        pipe_stage_90[0] = shift_reg[90] * COEFF_90;
        pipe_stage_91[0] = shift_reg[91] * COEFF_91;
        pipe_stage_92[0] = shift_reg[92] * COEFF_92;
        pipe_stage_93[0] = shift_reg[93] * COEFF_93;
        pipe_stage_94[0] = shift_reg[94] * COEFF_94;
        pipe_stage_95[0] = shift_reg[95] * COEFF_95;
        pipe_stage_96[0] = shift_reg[96] * COEFF_96;
        pipe_stage_97[0] = shift_reg[97] * COEFF_97;
        pipe_stage_98[0] = shift_reg[98] * COEFF_98;
        pipe_stage_99[0] = shift_reg[99] * COEFF_99;
        data_out = 0;
        data_out = data_out + pipe_stage_0[0];
        data_out = data_out + pipe_stage_1[0];
        data_out = data_out + pipe_stage_2[0];
        data_out = data_out + pipe_stage_3[0];
        data_out = data_out + pipe_stage_4[0];
        data_out = data_out + pipe_stage_5[0];
        data_out = data_out + pipe_stage_6[0];
        data_out = data_out + pipe_stage_7[0];
        data_out = data_out + pipe_stage_8[0];
        data_out = data_out + pipe_stage_9[0];
        data_out = data_out + pipe_stage_10[0];
        data_out = data_out + pipe_stage_11[0];
        data_out = data_out + pipe_stage_12[0];
        data_out = data_out + pipe_stage_13[0];
        data_out = data_out + pipe_stage_14[0];
        data_out = data_out + pipe_stage_15[0];
        data_out = data_out + pipe_stage_16[0];
        data_out = data_out + pipe_stage_17[0];
        data_out = data_out + pipe_stage_18[0];
        data_out = data_out + pipe_stage_19[0];
        data_out = data_out + pipe_stage_20[0];
        data_out = data_out + pipe_stage_21[0];
        data_out = data_out + pipe_stage_22[0];
        data_out = data_out + pipe_stage_23[0];
        data_out = data_out + pipe_stage_24[0];
        data_out = data_out + pipe_stage_25[0];
        data_out = data_out + pipe_stage_26[0];
        data_out = data_out + pipe_stage_27[0];
        data_out = data_out + pipe_stage_28[0];
        data_out = data_out + pipe_stage_29[0];
        data_out = data_out + pipe_stage_30[0];
        data_out = data_out + pipe_stage_31[0];
        data_out = data_out + pipe_stage_32[0];
        data_out = data_out + pipe_stage_33[0];
        data_out = data_out + pipe_stage_34[0];
        data_out = data_out + pipe_stage_35[0];
        data_out = data_out + pipe_stage_36[0];
        data_out = data_out + pipe_stage_37[0];
        data_out = data_out + pipe_stage_38[0];
        data_out = data_out + pipe_stage_39[0];
        data_out = data_out + pipe_stage_40[0];
        data_out = data_out + pipe_stage_41[0];
        data_out = data_out + pipe_stage_42[0];
        data_out = data_out + pipe_stage_43[0];
        data_out = data_out + pipe_stage_44[0];
        data_out = data_out + pipe_stage_45[0];
        data_out = data_out + pipe_stage_46[0];
        data_out = data_out + pipe_stage_47[0];
        data_out = data_out + pipe_stage_48[0];
        data_out = data_out + pipe_stage_49[0];
        data_out = data_out + pipe_stage_50[0];
        data_out = data_out + pipe_stage_51[0];
        data_out = data_out + pipe_stage_52[0];
        data_out = data_out + pipe_stage_53[0];
        data_out = data_out + pipe_stage_54[0];
        data_out = data_out + pipe_stage_55[0];
        data_out = data_out + pipe_stage_56[0];
        data_out = data_out + pipe_stage_57[0];
        data_out = data_out + pipe_stage_58[0];
        data_out = data_out + pipe_stage_59[0];
        data_out = data_out + pipe_stage_60[0];
        data_out = data_out + pipe_stage_61[0];
        data_out = data_out + pipe_stage_62[0];
        data_out = data_out + pipe_stage_63[0];
        data_out = data_out + pipe_stage_64[0];
        data_out = data_out + pipe_stage_65[0];
        data_out = data_out + pipe_stage_66[0];
        data_out = data_out + pipe_stage_67[0];
        data_out = data_out + pipe_stage_68[0];
        data_out = data_out + pipe_stage_69[0];
        data_out = data_out + pipe_stage_70[0];
        data_out = data_out + pipe_stage_71[0];
        data_out = data_out + pipe_stage_72[0];
        data_out = data_out + pipe_stage_73[0];
        data_out = data_out + pipe_stage_74[0];
        data_out = data_out + pipe_stage_75[0];
        data_out = data_out + pipe_stage_76[0];
        data_out = data_out + pipe_stage_77[0];
        data_out = data_out + pipe_stage_78[0];
        data_out = data_out + pipe_stage_79[0];
        data_out = data_out + pipe_stage_80[0];
        data_out = data_out + pipe_stage_81[0];
        data_out = data_out + pipe_stage_82[0];
        data_out = data_out + pipe_stage_83[0];
        data_out = data_out + pipe_stage_84[0];
        data_out = data_out + pipe_stage_85[0];
        data_out = data_out + pipe_stage_86[0];
        data_out = data_out + pipe_stage_87[0];
        data_out = data_out + pipe_stage_88[0];
        data_out = data_out + pipe_stage_89[0];
        data_out = data_out + pipe_stage_90[0];
        data_out = data_out + pipe_stage_91[0];
        data_out = data_out + pipe_stage_92[0];
        data_out = data_out + pipe_stage_93[0];
        data_out = data_out + pipe_stage_94[0];
        data_out = data_out + pipe_stage_95[0];
        data_out = data_out + pipe_stage_96[0];
        data_out = data_out + pipe_stage_97[0];
        data_out = data_out + pipe_stage_98[0];
        data_out = data_out + pipe_stage_99[0];

    end
end

endmodule
