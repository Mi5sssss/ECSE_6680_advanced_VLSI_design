
module fir_filter (
    input wire clk,                 // Clock signal
    input wire rst,                 // Reset signal
    input wire signed [15:0] data_in, // 16-bit signed input data
    output reg signed [31:0] data_out // 32-bit signed output data
);

// Number of taps
localparam TAPS = 336;
localparam signed [15:0] COEFF_0 = 16'sd0;
localparam signed [15:0] COEFF_1 = -16'sd0;
localparam signed [15:0] COEFF_2 = -16'sd0;
localparam signed [15:0] COEFF_3 = -16'sd0;
localparam signed [15:0] COEFF_4 = -16'sd0;
localparam signed [15:0] COEFF_5 = 16'sd0;
localparam signed [15:0] COEFF_6 = 16'sd0;
localparam signed [15:0] COEFF_7 = 16'sd0;
localparam signed [15:0] COEFF_8 = 16'sd0;
localparam signed [15:0] COEFF_9 = 16'sd0;
localparam signed [15:0] COEFF_10 = -16'sd0;
localparam signed [15:0] COEFF_11 = -16'sd0;
localparam signed [15:0] COEFF_12 = -16'sd0;
localparam signed [15:0] COEFF_13 = -16'sd0;
localparam signed [15:0] COEFF_14 = -16'sd0;
localparam signed [15:0] COEFF_15 = 16'sd0;
localparam signed [15:0] COEFF_16 = 16'sd1;
localparam signed [15:0] COEFF_17 = 16'sd1;
localparam signed [15:0] COEFF_18 = 16'sd0;
localparam signed [15:0] COEFF_19 = -16'sd0;
localparam signed [15:0] COEFF_20 = -16'sd1;
localparam signed [15:0] COEFF_21 = -16'sd1;
localparam signed [15:0] COEFF_22 = -16'sd1;
localparam signed [15:0] COEFF_23 = -16'sd0;
localparam signed [15:0] COEFF_24 = 16'sd1;
localparam signed [15:0] COEFF_25 = 16'sd2;
localparam signed [15:0] COEFF_26 = 16'sd2;
localparam signed [15:0] COEFF_27 = 16'sd1;
localparam signed [15:0] COEFF_28 = -16'sd0;
localparam signed [15:0] COEFF_29 = -16'sd2;
localparam signed [15:0] COEFF_30 = -16'sd3;
localparam signed [15:0] COEFF_31 = -16'sd3;
localparam signed [15:0] COEFF_32 = -16'sd1;
localparam signed [15:0] COEFF_33 = 16'sd1;
localparam signed [15:0] COEFF_34 = 16'sd3;
localparam signed [15:0] COEFF_35 = 16'sd4;
localparam signed [15:0] COEFF_36 = 16'sd3;
localparam signed [15:0] COEFF_37 = 16'sd0;
localparam signed [15:0] COEFF_38 = -16'sd2;
localparam signed [15:0] COEFF_39 = -16'sd5;
localparam signed [15:0] COEFF_40 = -16'sd6;
localparam signed [15:0] COEFF_41 = -16'sd3;
localparam signed [15:0] COEFF_42 = 16'sd0;
localparam signed [15:0] COEFF_43 = 16'sd5;
localparam signed [15:0] COEFF_44 = 16'sd7;
localparam signed [15:0] COEFF_45 = 16'sd7;
localparam signed [15:0] COEFF_46 = 16'sd3;
localparam signed [15:0] COEFF_47 = -16'sd2;
localparam signed [15:0] COEFF_48 = -16'sd8;
localparam signed [15:0] COEFF_49 = -16'sd10;
localparam signed [15:0] COEFF_50 = -16'sd8;
localparam signed [15:0] COEFF_51 = -16'sd1;
localparam signed [15:0] COEFF_52 = 16'sd6;
localparam signed [15:0] COEFF_53 = 16'sd11;
localparam signed [15:0] COEFF_54 = 16'sd12;
localparam signed [15:0] COEFF_55 = 16'sd7;
localparam signed [15:0] COEFF_56 = -16'sd1;
localparam signed [15:0] COEFF_57 = -16'sd10;
localparam signed [15:0] COEFF_58 = -16'sd16;
localparam signed [15:0] COEFF_59 = -16'sd14;
localparam signed [15:0] COEFF_60 = -16'sd6;
localparam signed [15:0] COEFF_61 = 16'sd5;
localparam signed [15:0] COEFF_62 = 16'sd16;
localparam signed [15:0] COEFF_63 = 16'sd20;
localparam signed [15:0] COEFF_64 = 16'sd15;
localparam signed [15:0] COEFF_65 = 16'sd2;
localparam signed [15:0] COEFF_66 = -16'sd12;
localparam signed [15:0] COEFF_67 = -16'sd22;
localparam signed [15:0] COEFF_68 = -16'sd23;
localparam signed [15:0] COEFF_69 = -16'sd13;
localparam signed [15:0] COEFF_70 = 16'sd3;
localparam signed [15:0] COEFF_71 = 16'sd20;
localparam signed [15:0] COEFF_72 = 16'sd29;
localparam signed [15:0] COEFF_73 = 16'sd26;
localparam signed [15:0] COEFF_74 = 16'sd10;
localparam signed [15:0] COEFF_75 = -16'sd11;
localparam signed [15:0] COEFF_76 = -16'sd29;
localparam signed [15:0] COEFF_77 = -16'sd35;
localparam signed [15:0] COEFF_78 = -16'sd26;
localparam signed [15:0] COEFF_79 = -16'sd3;
localparam signed [15:0] COEFF_80 = 16'sd22;
localparam signed [15:0] COEFF_81 = 16'sd40;
localparam signed [15:0] COEFF_82 = 16'sd40;
localparam signed [15:0] COEFF_83 = 16'sd22;
localparam signed [15:0] COEFF_84 = -16'sd7;
localparam signed [15:0] COEFF_85 = -16'sd36;
localparam signed [15:0] COEFF_86 = -16'sd50;
localparam signed [15:0] COEFF_87 = -16'sd43;
localparam signed [15:0] COEFF_88 = -16'sd15;
localparam signed [15:0] COEFF_89 = 16'sd21;
localparam signed [15:0] COEFF_90 = 16'sd51;
localparam signed [15:0] COEFF_91 = 16'sd60;
localparam signed [15:0] COEFF_92 = 16'sd42;
localparam signed [15:0] COEFF_93 = 16'sd3;
localparam signed [15:0] COEFF_94 = -16'sd39;
localparam signed [15:0] COEFF_95 = -16'sd67;
localparam signed [15:0] COEFF_96 = -16'sd66;
localparam signed [15:0] COEFF_97 = -16'sd35;
localparam signed [15:0] COEFF_98 = 16'sd13;
localparam signed [15:0] COEFF_99 = 16'sd60;
localparam signed [15:0] COEFF_100 = 16'sd83;
localparam signed [15:0] COEFF_101 = 16'sd69;
localparam signed [15:0] COEFF_102 = 16'sd22;
localparam signed [15:0] COEFF_103 = -16'sd37;
localparam signed [15:0] COEFF_104 = -16'sd84;
localparam signed [15:0] COEFF_105 = -16'sd96;
localparam signed [15:0] COEFF_106 = -16'sd65;
localparam signed [15:0] COEFF_107 = -16'sd2;
localparam signed [15:0] COEFF_108 = 16'sd65;
localparam signed [15:0] COEFF_109 = 16'sd109;
localparam signed [15:0] COEFF_110 = 16'sd105;
localparam signed [15:0] COEFF_111 = 16'sd53;
localparam signed [15:0] COEFF_112 = -16'sd26;
localparam signed [15:0] COEFF_113 = -16'sd99;
localparam signed [15:0] COEFF_114 = -16'sd132;
localparam signed [15:0] COEFF_115 = -16'sd107;
localparam signed [15:0] COEFF_116 = -16'sd32;
localparam signed [15:0] COEFF_117 = 16'sd63;
localparam signed [15:0] COEFF_118 = 16'sd136;
localparam signed [15:0] COEFF_119 = 16'sd153;
localparam signed [15:0] COEFF_120 = 16'sd100;
localparam signed [15:0] COEFF_121 = -16'sd1;
localparam signed [15:0] COEFF_122 = -16'sd109;
localparam signed [15:0] COEFF_123 = -16'sd176;
localparam signed [15:0] COEFF_124 = -16'sd166;
localparam signed [15:0] COEFF_125 = -16'sd80;
localparam signed [15:0] COEFF_126 = 16'sd48;
localparam signed [15:0] COEFF_127 = 16'sd164;
localparam signed [15:0] COEFF_128 = 16'sd214;
localparam signed [15:0] COEFF_129 = 16'sd170;
localparam signed [15:0] COEFF_130 = 16'sd45;
localparam signed [15:0] COEFF_131 = -16'sd110;
localparam signed [15:0] COEFF_132 = -16'sd227;
localparam signed [15:0] COEFF_133 = -16'sd249;
localparam signed [15:0] COEFF_134 = -16'sd159;
localparam signed [15:0] COEFF_135 = 16'sd10;
localparam signed [15:0] COEFF_136 = 16'sd190;
localparam signed [15:0] COEFF_137 = 16'sd297;
localparam signed [15:0] COEFF_138 = 16'sd277;
localparam signed [15:0] COEFF_139 = 16'sd128;
localparam signed [15:0] COEFF_140 = -16'sd93;
localparam signed [15:0] COEFF_141 = -16'sd291;
localparam signed [15:0] COEFF_142 = -16'sd374;
localparam signed [15:0] COEFF_143 = -16'sd293;
localparam signed [15:0] COEFF_144 = -16'sd67;
localparam signed [15:0] COEFF_145 = 16'sd211;
localparam signed [15:0] COEFF_146 = 16'sd423;
localparam signed [15:0] COEFF_147 = 16'sd461;
localparam signed [15:0] COEFF_148 = 16'sd289;
localparam signed [15:0] COEFF_149 = -16'sd38;
localparam signed [15:0] COEFF_150 = -16'sd388;
localparam signed [15:0] COEFF_151 = -16'sd603;
localparam signed [15:0] COEFF_152 = -16'sd563;
localparam signed [15:0] COEFF_153 = -16'sd252;
localparam signed [15:0] COEFF_154 = 16'sd227;
localparam signed [15:0] COEFF_155 = 16'sd679;
localparam signed [15:0] COEFF_156 = 16'sd888;
localparam signed [15:0] COEFF_157 = 16'sd708;
localparam signed [15:0] COEFF_158 = 16'sd144;
localparam signed [15:0] COEFF_159 = -16'sd626;
localparam signed [15:0] COEFF_160 = -16'sd1295;
localparam signed [15:0] COEFF_161 = -16'sd1513;
localparam signed [15:0] COEFF_162 = -16'sd1024;
localparam signed [15:0] COEFF_163 = 16'sd235;
localparam signed [15:0] COEFF_164 = 16'sd2087;
localparam signed [15:0] COEFF_165 = 16'sd4139;
localparam signed [15:0] COEFF_166 = 16'sd5898;
localparam signed [15:0] COEFF_167 = 16'sd6911;
localparam signed [15:0] COEFF_168 = 16'sd6911;
localparam signed [15:0] COEFF_169 = 16'sd5898;
localparam signed [15:0] COEFF_170 = 16'sd4139;
localparam signed [15:0] COEFF_171 = 16'sd2087;
localparam signed [15:0] COEFF_172 = 16'sd235;
localparam signed [15:0] COEFF_173 = -16'sd1024;
localparam signed [15:0] COEFF_174 = -16'sd1513;
localparam signed [15:0] COEFF_175 = -16'sd1295;
localparam signed [15:0] COEFF_176 = -16'sd626;
localparam signed [15:0] COEFF_177 = 16'sd144;
localparam signed [15:0] COEFF_178 = 16'sd708;
localparam signed [15:0] COEFF_179 = 16'sd888;
localparam signed [15:0] COEFF_180 = 16'sd679;
localparam signed [15:0] COEFF_181 = 16'sd227;
localparam signed [15:0] COEFF_182 = -16'sd252;
localparam signed [15:0] COEFF_183 = -16'sd563;
localparam signed [15:0] COEFF_184 = -16'sd603;
localparam signed [15:0] COEFF_185 = -16'sd388;
localparam signed [15:0] COEFF_186 = -16'sd38;
localparam signed [15:0] COEFF_187 = 16'sd289;
localparam signed [15:0] COEFF_188 = 16'sd461;
localparam signed [15:0] COEFF_189 = 16'sd423;
localparam signed [15:0] COEFF_190 = 16'sd211;
localparam signed [15:0] COEFF_191 = -16'sd67;
localparam signed [15:0] COEFF_192 = -16'sd293;
localparam signed [15:0] COEFF_193 = -16'sd374;
localparam signed [15:0] COEFF_194 = -16'sd291;
localparam signed [15:0] COEFF_195 = -16'sd93;
localparam signed [15:0] COEFF_196 = 16'sd128;
localparam signed [15:0] COEFF_197 = 16'sd277;
localparam signed [15:0] COEFF_198 = 16'sd297;
localparam signed [15:0] COEFF_199 = 16'sd190;
localparam signed [15:0] COEFF_200 = 16'sd10;
localparam signed [15:0] COEFF_201 = -16'sd159;
localparam signed [15:0] COEFF_202 = -16'sd249;
localparam signed [15:0] COEFF_203 = -16'sd227;
localparam signed [15:0] COEFF_204 = -16'sd110;
localparam signed [15:0] COEFF_205 = 16'sd45;
localparam signed [15:0] COEFF_206 = 16'sd170;
localparam signed [15:0] COEFF_207 = 16'sd214;
localparam signed [15:0] COEFF_208 = 16'sd164;
localparam signed [15:0] COEFF_209 = 16'sd48;
localparam signed [15:0] COEFF_210 = -16'sd80;
localparam signed [15:0] COEFF_211 = -16'sd166;
localparam signed [15:0] COEFF_212 = -16'sd176;
localparam signed [15:0] COEFF_213 = -16'sd109;
localparam signed [15:0] COEFF_214 = -16'sd1;
localparam signed [15:0] COEFF_215 = 16'sd100;
localparam signed [15:0] COEFF_216 = 16'sd153;
localparam signed [15:0] COEFF_217 = 16'sd136;
localparam signed [15:0] COEFF_218 = 16'sd63;
localparam signed [15:0] COEFF_219 = -16'sd32;
localparam signed [15:0] COEFF_220 = -16'sd107;
localparam signed [15:0] COEFF_221 = -16'sd132;
localparam signed [15:0] COEFF_222 = -16'sd99;
localparam signed [15:0] COEFF_223 = -16'sd26;
localparam signed [15:0] COEFF_224 = 16'sd53;
localparam signed [15:0] COEFF_225 = 16'sd105;
localparam signed [15:0] COEFF_226 = 16'sd109;
localparam signed [15:0] COEFF_227 = 16'sd65;
localparam signed [15:0] COEFF_228 = -16'sd2;
localparam signed [15:0] COEFF_229 = -16'sd65;
localparam signed [15:0] COEFF_230 = -16'sd96;
localparam signed [15:0] COEFF_231 = -16'sd84;
localparam signed [15:0] COEFF_232 = -16'sd37;
localparam signed [15:0] COEFF_233 = 16'sd22;
localparam signed [15:0] COEFF_234 = 16'sd69;
localparam signed [15:0] COEFF_235 = 16'sd83;
localparam signed [15:0] COEFF_236 = 16'sd60;
localparam signed [15:0] COEFF_237 = 16'sd13;
localparam signed [15:0] COEFF_238 = -16'sd35;
localparam signed [15:0] COEFF_239 = -16'sd66;
localparam signed [15:0] COEFF_240 = -16'sd67;
localparam signed [15:0] COEFF_241 = -16'sd39;
localparam signed [15:0] COEFF_242 = 16'sd3;
localparam signed [15:0] COEFF_243 = 16'sd42;
localparam signed [15:0] COEFF_244 = 16'sd60;
localparam signed [15:0] COEFF_245 = 16'sd51;
localparam signed [15:0] COEFF_246 = 16'sd21;
localparam signed [15:0] COEFF_247 = -16'sd15;
localparam signed [15:0] COEFF_248 = -16'sd43;
localparam signed [15:0] COEFF_249 = -16'sd50;
localparam signed [15:0] COEFF_250 = -16'sd36;
localparam signed [15:0] COEFF_251 = -16'sd7;
localparam signed [15:0] COEFF_252 = 16'sd22;
localparam signed [15:0] COEFF_253 = 16'sd40;
localparam signed [15:0] COEFF_254 = 16'sd40;
localparam signed [15:0] COEFF_255 = 16'sd22;
localparam signed [15:0] COEFF_256 = -16'sd3;
localparam signed [15:0] COEFF_257 = -16'sd26;
localparam signed [15:0] COEFF_258 = -16'sd35;
localparam signed [15:0] COEFF_259 = -16'sd29;
localparam signed [15:0] COEFF_260 = -16'sd11;
localparam signed [15:0] COEFF_261 = 16'sd10;
localparam signed [15:0] COEFF_262 = 16'sd26;
localparam signed [15:0] COEFF_263 = 16'sd29;
localparam signed [15:0] COEFF_264 = 16'sd20;
localparam signed [15:0] COEFF_265 = 16'sd3;
localparam signed [15:0] COEFF_266 = -16'sd13;
localparam signed [15:0] COEFF_267 = -16'sd23;
localparam signed [15:0] COEFF_268 = -16'sd22;
localparam signed [15:0] COEFF_269 = -16'sd12;
localparam signed [15:0] COEFF_270 = 16'sd2;
localparam signed [15:0] COEFF_271 = 16'sd15;
localparam signed [15:0] COEFF_272 = 16'sd20;
localparam signed [15:0] COEFF_273 = 16'sd16;
localparam signed [15:0] COEFF_274 = 16'sd5;
localparam signed [15:0] COEFF_275 = -16'sd6;
localparam signed [15:0] COEFF_276 = -16'sd14;
localparam signed [15:0] COEFF_277 = -16'sd16;
localparam signed [15:0] COEFF_278 = -16'sd10;
localparam signed [15:0] COEFF_279 = -16'sd1;
localparam signed [15:0] COEFF_280 = 16'sd7;
localparam signed [15:0] COEFF_281 = 16'sd12;
localparam signed [15:0] COEFF_282 = 16'sd11;
localparam signed [15:0] COEFF_283 = 16'sd6;
localparam signed [15:0] COEFF_284 = -16'sd1;
localparam signed [15:0] COEFF_285 = -16'sd8;
localparam signed [15:0] COEFF_286 = -16'sd10;
localparam signed [15:0] COEFF_287 = -16'sd8;
localparam signed [15:0] COEFF_288 = -16'sd2;
localparam signed [15:0] COEFF_289 = 16'sd3;
localparam signed [15:0] COEFF_290 = 16'sd7;
localparam signed [15:0] COEFF_291 = 16'sd7;
localparam signed [15:0] COEFF_292 = 16'sd5;
localparam signed [15:0] COEFF_293 = 16'sd0;
localparam signed [15:0] COEFF_294 = -16'sd3;
localparam signed [15:0] COEFF_295 = -16'sd6;
localparam signed [15:0] COEFF_296 = -16'sd5;
localparam signed [15:0] COEFF_297 = -16'sd2;
localparam signed [15:0] COEFF_298 = 16'sd0;
localparam signed [15:0] COEFF_299 = 16'sd3;
localparam signed [15:0] COEFF_300 = 16'sd4;
localparam signed [15:0] COEFF_301 = 16'sd3;
localparam signed [15:0] COEFF_302 = 16'sd1;
localparam signed [15:0] COEFF_303 = -16'sd1;
localparam signed [15:0] COEFF_304 = -16'sd3;
localparam signed [15:0] COEFF_305 = -16'sd3;
localparam signed [15:0] COEFF_306 = -16'sd2;
localparam signed [15:0] COEFF_307 = -16'sd0;
localparam signed [15:0] COEFF_308 = 16'sd1;
localparam signed [15:0] COEFF_309 = 16'sd2;
localparam signed [15:0] COEFF_310 = 16'sd2;
localparam signed [15:0] COEFF_311 = 16'sd1;
localparam signed [15:0] COEFF_312 = -16'sd0;
localparam signed [15:0] COEFF_313 = -16'sd1;
localparam signed [15:0] COEFF_314 = -16'sd1;
localparam signed [15:0] COEFF_315 = -16'sd1;
localparam signed [15:0] COEFF_316 = -16'sd0;
localparam signed [15:0] COEFF_317 = 16'sd0;
localparam signed [15:0] COEFF_318 = 16'sd1;
localparam signed [15:0] COEFF_319 = 16'sd1;
localparam signed [15:0] COEFF_320 = 16'sd0;
localparam signed [15:0] COEFF_321 = -16'sd0;
localparam signed [15:0] COEFF_322 = -16'sd0;
localparam signed [15:0] COEFF_323 = -16'sd0;
localparam signed [15:0] COEFF_324 = -16'sd0;
localparam signed [15:0] COEFF_325 = -16'sd0;
localparam signed [15:0] COEFF_326 = 16'sd0;
localparam signed [15:0] COEFF_327 = 16'sd0;
localparam signed [15:0] COEFF_328 = 16'sd0;
localparam signed [15:0] COEFF_329 = 16'sd0;
localparam signed [15:0] COEFF_330 = 16'sd0;
localparam signed [15:0] COEFF_331 = -16'sd0;
localparam signed [15:0] COEFF_332 = -16'sd0;
localparam signed [15:0] COEFF_333 = -16'sd0;
localparam signed [15:0] COEFF_334 = -16'sd0;
localparam signed [15:0] COEFF_335 = 16'sd0;

// Shift register for input samples
reg signed [15:0] shift_reg[TAPS-1:0];
reg signed [31:0] temp_data_out;  // Temporary variable for accumulation

// Multiply and accumulate
integer i;
always @(posedge clk) begin
    if (rst) begin
        // Clear the shift register and temporary accumulator
        for (i = 0; i < TAPS; i = i + 1) begin
            shift_reg[i] <= 0;
        end
        temp_data_out <= 0;
        data_out <= 0;
    end else begin
        // Shift the input sample through the register
        for (i = TAPS-1; i > 0; i = i - 1) begin
            shift_reg[i] <= shift_reg[i - 1];
        end
        shift_reg[0] <= data_in;

        // Initialize the accumulator at the start of each cycle
        temp_data_out = 0;
        temp_data_out = temp_data_out + shift_reg[0] * COEFF_0;
        temp_data_out = temp_data_out + shift_reg[1] * COEFF_1;
        temp_data_out = temp_data_out + shift_reg[2] * COEFF_2;
        temp_data_out = temp_data_out + shift_reg[3] * COEFF_3;
        temp_data_out = temp_data_out + shift_reg[4] * COEFF_4;
        temp_data_out = temp_data_out + shift_reg[5] * COEFF_5;
        temp_data_out = temp_data_out + shift_reg[6] * COEFF_6;
        temp_data_out = temp_data_out + shift_reg[7] * COEFF_7;
        temp_data_out = temp_data_out + shift_reg[8] * COEFF_8;
        temp_data_out = temp_data_out + shift_reg[9] * COEFF_9;
        temp_data_out = temp_data_out + shift_reg[10] * COEFF_10;
        temp_data_out = temp_data_out + shift_reg[11] * COEFF_11;
        temp_data_out = temp_data_out + shift_reg[12] * COEFF_12;
        temp_data_out = temp_data_out + shift_reg[13] * COEFF_13;
        temp_data_out = temp_data_out + shift_reg[14] * COEFF_14;
        temp_data_out = temp_data_out + shift_reg[15] * COEFF_15;
        temp_data_out = temp_data_out + shift_reg[16] * COEFF_16;
        temp_data_out = temp_data_out + shift_reg[17] * COEFF_17;
        temp_data_out = temp_data_out + shift_reg[18] * COEFF_18;
        temp_data_out = temp_data_out + shift_reg[19] * COEFF_19;
        temp_data_out = temp_data_out + shift_reg[20] * COEFF_20;
        temp_data_out = temp_data_out + shift_reg[21] * COEFF_21;
        temp_data_out = temp_data_out + shift_reg[22] * COEFF_22;
        temp_data_out = temp_data_out + shift_reg[23] * COEFF_23;
        temp_data_out = temp_data_out + shift_reg[24] * COEFF_24;
        temp_data_out = temp_data_out + shift_reg[25] * COEFF_25;
        temp_data_out = temp_data_out + shift_reg[26] * COEFF_26;
        temp_data_out = temp_data_out + shift_reg[27] * COEFF_27;
        temp_data_out = temp_data_out + shift_reg[28] * COEFF_28;
        temp_data_out = temp_data_out + shift_reg[29] * COEFF_29;
        temp_data_out = temp_data_out + shift_reg[30] * COEFF_30;
        temp_data_out = temp_data_out + shift_reg[31] * COEFF_31;
        temp_data_out = temp_data_out + shift_reg[32] * COEFF_32;
        temp_data_out = temp_data_out + shift_reg[33] * COEFF_33;
        temp_data_out = temp_data_out + shift_reg[34] * COEFF_34;
        temp_data_out = temp_data_out + shift_reg[35] * COEFF_35;
        temp_data_out = temp_data_out + shift_reg[36] * COEFF_36;
        temp_data_out = temp_data_out + shift_reg[37] * COEFF_37;
        temp_data_out = temp_data_out + shift_reg[38] * COEFF_38;
        temp_data_out = temp_data_out + shift_reg[39] * COEFF_39;
        temp_data_out = temp_data_out + shift_reg[40] * COEFF_40;
        temp_data_out = temp_data_out + shift_reg[41] * COEFF_41;
        temp_data_out = temp_data_out + shift_reg[42] * COEFF_42;
        temp_data_out = temp_data_out + shift_reg[43] * COEFF_43;
        temp_data_out = temp_data_out + shift_reg[44] * COEFF_44;
        temp_data_out = temp_data_out + shift_reg[45] * COEFF_45;
        temp_data_out = temp_data_out + shift_reg[46] * COEFF_46;
        temp_data_out = temp_data_out + shift_reg[47] * COEFF_47;
        temp_data_out = temp_data_out + shift_reg[48] * COEFF_48;
        temp_data_out = temp_data_out + shift_reg[49] * COEFF_49;
        temp_data_out = temp_data_out + shift_reg[50] * COEFF_50;
        temp_data_out = temp_data_out + shift_reg[51] * COEFF_51;
        temp_data_out = temp_data_out + shift_reg[52] * COEFF_52;
        temp_data_out = temp_data_out + shift_reg[53] * COEFF_53;
        temp_data_out = temp_data_out + shift_reg[54] * COEFF_54;
        temp_data_out = temp_data_out + shift_reg[55] * COEFF_55;
        temp_data_out = temp_data_out + shift_reg[56] * COEFF_56;
        temp_data_out = temp_data_out + shift_reg[57] * COEFF_57;
        temp_data_out = temp_data_out + shift_reg[58] * COEFF_58;
        temp_data_out = temp_data_out + shift_reg[59] * COEFF_59;
        temp_data_out = temp_data_out + shift_reg[60] * COEFF_60;
        temp_data_out = temp_data_out + shift_reg[61] * COEFF_61;
        temp_data_out = temp_data_out + shift_reg[62] * COEFF_62;
        temp_data_out = temp_data_out + shift_reg[63] * COEFF_63;
        temp_data_out = temp_data_out + shift_reg[64] * COEFF_64;
        temp_data_out = temp_data_out + shift_reg[65] * COEFF_65;
        temp_data_out = temp_data_out + shift_reg[66] * COEFF_66;
        temp_data_out = temp_data_out + shift_reg[67] * COEFF_67;
        temp_data_out = temp_data_out + shift_reg[68] * COEFF_68;
        temp_data_out = temp_data_out + shift_reg[69] * COEFF_69;
        temp_data_out = temp_data_out + shift_reg[70] * COEFF_70;
        temp_data_out = temp_data_out + shift_reg[71] * COEFF_71;
        temp_data_out = temp_data_out + shift_reg[72] * COEFF_72;
        temp_data_out = temp_data_out + shift_reg[73] * COEFF_73;
        temp_data_out = temp_data_out + shift_reg[74] * COEFF_74;
        temp_data_out = temp_data_out + shift_reg[75] * COEFF_75;
        temp_data_out = temp_data_out + shift_reg[76] * COEFF_76;
        temp_data_out = temp_data_out + shift_reg[77] * COEFF_77;
        temp_data_out = temp_data_out + shift_reg[78] * COEFF_78;
        temp_data_out = temp_data_out + shift_reg[79] * COEFF_79;
        temp_data_out = temp_data_out + shift_reg[80] * COEFF_80;
        temp_data_out = temp_data_out + shift_reg[81] * COEFF_81;
        temp_data_out = temp_data_out + shift_reg[82] * COEFF_82;
        temp_data_out = temp_data_out + shift_reg[83] * COEFF_83;
        temp_data_out = temp_data_out + shift_reg[84] * COEFF_84;
        temp_data_out = temp_data_out + shift_reg[85] * COEFF_85;
        temp_data_out = temp_data_out + shift_reg[86] * COEFF_86;
        temp_data_out = temp_data_out + shift_reg[87] * COEFF_87;
        temp_data_out = temp_data_out + shift_reg[88] * COEFF_88;
        temp_data_out = temp_data_out + shift_reg[89] * COEFF_89;
        temp_data_out = temp_data_out + shift_reg[90] * COEFF_90;
        temp_data_out = temp_data_out + shift_reg[91] * COEFF_91;
        temp_data_out = temp_data_out + shift_reg[92] * COEFF_92;
        temp_data_out = temp_data_out + shift_reg[93] * COEFF_93;
        temp_data_out = temp_data_out + shift_reg[94] * COEFF_94;
        temp_data_out = temp_data_out + shift_reg[95] * COEFF_95;
        temp_data_out = temp_data_out + shift_reg[96] * COEFF_96;
        temp_data_out = temp_data_out + shift_reg[97] * COEFF_97;
        temp_data_out = temp_data_out + shift_reg[98] * COEFF_98;
        temp_data_out = temp_data_out + shift_reg[99] * COEFF_99;
        temp_data_out = temp_data_out + shift_reg[100] * COEFF_100;
        temp_data_out = temp_data_out + shift_reg[101] * COEFF_101;
        temp_data_out = temp_data_out + shift_reg[102] * COEFF_102;
        temp_data_out = temp_data_out + shift_reg[103] * COEFF_103;
        temp_data_out = temp_data_out + shift_reg[104] * COEFF_104;
        temp_data_out = temp_data_out + shift_reg[105] * COEFF_105;
        temp_data_out = temp_data_out + shift_reg[106] * COEFF_106;
        temp_data_out = temp_data_out + shift_reg[107] * COEFF_107;
        temp_data_out = temp_data_out + shift_reg[108] * COEFF_108;
        temp_data_out = temp_data_out + shift_reg[109] * COEFF_109;
        temp_data_out = temp_data_out + shift_reg[110] * COEFF_110;
        temp_data_out = temp_data_out + shift_reg[111] * COEFF_111;
        temp_data_out = temp_data_out + shift_reg[112] * COEFF_112;
        temp_data_out = temp_data_out + shift_reg[113] * COEFF_113;
        temp_data_out = temp_data_out + shift_reg[114] * COEFF_114;
        temp_data_out = temp_data_out + shift_reg[115] * COEFF_115;
        temp_data_out = temp_data_out + shift_reg[116] * COEFF_116;
        temp_data_out = temp_data_out + shift_reg[117] * COEFF_117;
        temp_data_out = temp_data_out + shift_reg[118] * COEFF_118;
        temp_data_out = temp_data_out + shift_reg[119] * COEFF_119;
        temp_data_out = temp_data_out + shift_reg[120] * COEFF_120;
        temp_data_out = temp_data_out + shift_reg[121] * COEFF_121;
        temp_data_out = temp_data_out + shift_reg[122] * COEFF_122;
        temp_data_out = temp_data_out + shift_reg[123] * COEFF_123;
        temp_data_out = temp_data_out + shift_reg[124] * COEFF_124;
        temp_data_out = temp_data_out + shift_reg[125] * COEFF_125;
        temp_data_out = temp_data_out + shift_reg[126] * COEFF_126;
        temp_data_out = temp_data_out + shift_reg[127] * COEFF_127;
        temp_data_out = temp_data_out + shift_reg[128] * COEFF_128;
        temp_data_out = temp_data_out + shift_reg[129] * COEFF_129;
        temp_data_out = temp_data_out + shift_reg[130] * COEFF_130;
        temp_data_out = temp_data_out + shift_reg[131] * COEFF_131;
        temp_data_out = temp_data_out + shift_reg[132] * COEFF_132;
        temp_data_out = temp_data_out + shift_reg[133] * COEFF_133;
        temp_data_out = temp_data_out + shift_reg[134] * COEFF_134;
        temp_data_out = temp_data_out + shift_reg[135] * COEFF_135;
        temp_data_out = temp_data_out + shift_reg[136] * COEFF_136;
        temp_data_out = temp_data_out + shift_reg[137] * COEFF_137;
        temp_data_out = temp_data_out + shift_reg[138] * COEFF_138;
        temp_data_out = temp_data_out + shift_reg[139] * COEFF_139;
        temp_data_out = temp_data_out + shift_reg[140] * COEFF_140;
        temp_data_out = temp_data_out + shift_reg[141] * COEFF_141;
        temp_data_out = temp_data_out + shift_reg[142] * COEFF_142;
        temp_data_out = temp_data_out + shift_reg[143] * COEFF_143;
        temp_data_out = temp_data_out + shift_reg[144] * COEFF_144;
        temp_data_out = temp_data_out + shift_reg[145] * COEFF_145;
        temp_data_out = temp_data_out + shift_reg[146] * COEFF_146;
        temp_data_out = temp_data_out + shift_reg[147] * COEFF_147;
        temp_data_out = temp_data_out + shift_reg[148] * COEFF_148;
        temp_data_out = temp_data_out + shift_reg[149] * COEFF_149;
        temp_data_out = temp_data_out + shift_reg[150] * COEFF_150;
        temp_data_out = temp_data_out + shift_reg[151] * COEFF_151;
        temp_data_out = temp_data_out + shift_reg[152] * COEFF_152;
        temp_data_out = temp_data_out + shift_reg[153] * COEFF_153;
        temp_data_out = temp_data_out + shift_reg[154] * COEFF_154;
        temp_data_out = temp_data_out + shift_reg[155] * COEFF_155;
        temp_data_out = temp_data_out + shift_reg[156] * COEFF_156;
        temp_data_out = temp_data_out + shift_reg[157] * COEFF_157;
        temp_data_out = temp_data_out + shift_reg[158] * COEFF_158;
        temp_data_out = temp_data_out + shift_reg[159] * COEFF_159;
        temp_data_out = temp_data_out + shift_reg[160] * COEFF_160;
        temp_data_out = temp_data_out + shift_reg[161] * COEFF_161;
        temp_data_out = temp_data_out + shift_reg[162] * COEFF_162;
        temp_data_out = temp_data_out + shift_reg[163] * COEFF_163;
        temp_data_out = temp_data_out + shift_reg[164] * COEFF_164;
        temp_data_out = temp_data_out + shift_reg[165] * COEFF_165;
        temp_data_out = temp_data_out + shift_reg[166] * COEFF_166;
        temp_data_out = temp_data_out + shift_reg[167] * COEFF_167;
        temp_data_out = temp_data_out + shift_reg[168] * COEFF_168;
        temp_data_out = temp_data_out + shift_reg[169] * COEFF_169;
        temp_data_out = temp_data_out + shift_reg[170] * COEFF_170;
        temp_data_out = temp_data_out + shift_reg[171] * COEFF_171;
        temp_data_out = temp_data_out + shift_reg[172] * COEFF_172;
        temp_data_out = temp_data_out + shift_reg[173] * COEFF_173;
        temp_data_out = temp_data_out + shift_reg[174] * COEFF_174;
        temp_data_out = temp_data_out + shift_reg[175] * COEFF_175;
        temp_data_out = temp_data_out + shift_reg[176] * COEFF_176;
        temp_data_out = temp_data_out + shift_reg[177] * COEFF_177;
        temp_data_out = temp_data_out + shift_reg[178] * COEFF_178;
        temp_data_out = temp_data_out + shift_reg[179] * COEFF_179;
        temp_data_out = temp_data_out + shift_reg[180] * COEFF_180;
        temp_data_out = temp_data_out + shift_reg[181] * COEFF_181;
        temp_data_out = temp_data_out + shift_reg[182] * COEFF_182;
        temp_data_out = temp_data_out + shift_reg[183] * COEFF_183;
        temp_data_out = temp_data_out + shift_reg[184] * COEFF_184;
        temp_data_out = temp_data_out + shift_reg[185] * COEFF_185;
        temp_data_out = temp_data_out + shift_reg[186] * COEFF_186;
        temp_data_out = temp_data_out + shift_reg[187] * COEFF_187;
        temp_data_out = temp_data_out + shift_reg[188] * COEFF_188;
        temp_data_out = temp_data_out + shift_reg[189] * COEFF_189;
        temp_data_out = temp_data_out + shift_reg[190] * COEFF_190;
        temp_data_out = temp_data_out + shift_reg[191] * COEFF_191;
        temp_data_out = temp_data_out + shift_reg[192] * COEFF_192;
        temp_data_out = temp_data_out + shift_reg[193] * COEFF_193;
        temp_data_out = temp_data_out + shift_reg[194] * COEFF_194;
        temp_data_out = temp_data_out + shift_reg[195] * COEFF_195;
        temp_data_out = temp_data_out + shift_reg[196] * COEFF_196;
        temp_data_out = temp_data_out + shift_reg[197] * COEFF_197;
        temp_data_out = temp_data_out + shift_reg[198] * COEFF_198;
        temp_data_out = temp_data_out + shift_reg[199] * COEFF_199;
        temp_data_out = temp_data_out + shift_reg[200] * COEFF_200;
        temp_data_out = temp_data_out + shift_reg[201] * COEFF_201;
        temp_data_out = temp_data_out + shift_reg[202] * COEFF_202;
        temp_data_out = temp_data_out + shift_reg[203] * COEFF_203;
        temp_data_out = temp_data_out + shift_reg[204] * COEFF_204;
        temp_data_out = temp_data_out + shift_reg[205] * COEFF_205;
        temp_data_out = temp_data_out + shift_reg[206] * COEFF_206;
        temp_data_out = temp_data_out + shift_reg[207] * COEFF_207;
        temp_data_out = temp_data_out + shift_reg[208] * COEFF_208;
        temp_data_out = temp_data_out + shift_reg[209] * COEFF_209;
        temp_data_out = temp_data_out + shift_reg[210] * COEFF_210;
        temp_data_out = temp_data_out + shift_reg[211] * COEFF_211;
        temp_data_out = temp_data_out + shift_reg[212] * COEFF_212;
        temp_data_out = temp_data_out + shift_reg[213] * COEFF_213;
        temp_data_out = temp_data_out + shift_reg[214] * COEFF_214;
        temp_data_out = temp_data_out + shift_reg[215] * COEFF_215;
        temp_data_out = temp_data_out + shift_reg[216] * COEFF_216;
        temp_data_out = temp_data_out + shift_reg[217] * COEFF_217;
        temp_data_out = temp_data_out + shift_reg[218] * COEFF_218;
        temp_data_out = temp_data_out + shift_reg[219] * COEFF_219;
        temp_data_out = temp_data_out + shift_reg[220] * COEFF_220;
        temp_data_out = temp_data_out + shift_reg[221] * COEFF_221;
        temp_data_out = temp_data_out + shift_reg[222] * COEFF_222;
        temp_data_out = temp_data_out + shift_reg[223] * COEFF_223;
        temp_data_out = temp_data_out + shift_reg[224] * COEFF_224;
        temp_data_out = temp_data_out + shift_reg[225] * COEFF_225;
        temp_data_out = temp_data_out + shift_reg[226] * COEFF_226;
        temp_data_out = temp_data_out + shift_reg[227] * COEFF_227;
        temp_data_out = temp_data_out + shift_reg[228] * COEFF_228;
        temp_data_out = temp_data_out + shift_reg[229] * COEFF_229;
        temp_data_out = temp_data_out + shift_reg[230] * COEFF_230;
        temp_data_out = temp_data_out + shift_reg[231] * COEFF_231;
        temp_data_out = temp_data_out + shift_reg[232] * COEFF_232;
        temp_data_out = temp_data_out + shift_reg[233] * COEFF_233;
        temp_data_out = temp_data_out + shift_reg[234] * COEFF_234;
        temp_data_out = temp_data_out + shift_reg[235] * COEFF_235;
        temp_data_out = temp_data_out + shift_reg[236] * COEFF_236;
        temp_data_out = temp_data_out + shift_reg[237] * COEFF_237;
        temp_data_out = temp_data_out + shift_reg[238] * COEFF_238;
        temp_data_out = temp_data_out + shift_reg[239] * COEFF_239;
        temp_data_out = temp_data_out + shift_reg[240] * COEFF_240;
        temp_data_out = temp_data_out + shift_reg[241] * COEFF_241;
        temp_data_out = temp_data_out + shift_reg[242] * COEFF_242;
        temp_data_out = temp_data_out + shift_reg[243] * COEFF_243;
        temp_data_out = temp_data_out + shift_reg[244] * COEFF_244;
        temp_data_out = temp_data_out + shift_reg[245] * COEFF_245;
        temp_data_out = temp_data_out + shift_reg[246] * COEFF_246;
        temp_data_out = temp_data_out + shift_reg[247] * COEFF_247;
        temp_data_out = temp_data_out + shift_reg[248] * COEFF_248;
        temp_data_out = temp_data_out + shift_reg[249] * COEFF_249;
        temp_data_out = temp_data_out + shift_reg[250] * COEFF_250;
        temp_data_out = temp_data_out + shift_reg[251] * COEFF_251;
        temp_data_out = temp_data_out + shift_reg[252] * COEFF_252;
        temp_data_out = temp_data_out + shift_reg[253] * COEFF_253;
        temp_data_out = temp_data_out + shift_reg[254] * COEFF_254;
        temp_data_out = temp_data_out + shift_reg[255] * COEFF_255;
        temp_data_out = temp_data_out + shift_reg[256] * COEFF_256;
        temp_data_out = temp_data_out + shift_reg[257] * COEFF_257;
        temp_data_out = temp_data_out + shift_reg[258] * COEFF_258;
        temp_data_out = temp_data_out + shift_reg[259] * COEFF_259;
        temp_data_out = temp_data_out + shift_reg[260] * COEFF_260;
        temp_data_out = temp_data_out + shift_reg[261] * COEFF_261;
        temp_data_out = temp_data_out + shift_reg[262] * COEFF_262;
        temp_data_out = temp_data_out + shift_reg[263] * COEFF_263;
        temp_data_out = temp_data_out + shift_reg[264] * COEFF_264;
        temp_data_out = temp_data_out + shift_reg[265] * COEFF_265;
        temp_data_out = temp_data_out + shift_reg[266] * COEFF_266;
        temp_data_out = temp_data_out + shift_reg[267] * COEFF_267;
        temp_data_out = temp_data_out + shift_reg[268] * COEFF_268;
        temp_data_out = temp_data_out + shift_reg[269] * COEFF_269;
        temp_data_out = temp_data_out + shift_reg[270] * COEFF_270;
        temp_data_out = temp_data_out + shift_reg[271] * COEFF_271;
        temp_data_out = temp_data_out + shift_reg[272] * COEFF_272;
        temp_data_out = temp_data_out + shift_reg[273] * COEFF_273;
        temp_data_out = temp_data_out + shift_reg[274] * COEFF_274;
        temp_data_out = temp_data_out + shift_reg[275] * COEFF_275;
        temp_data_out = temp_data_out + shift_reg[276] * COEFF_276;
        temp_data_out = temp_data_out + shift_reg[277] * COEFF_277;
        temp_data_out = temp_data_out + shift_reg[278] * COEFF_278;
        temp_data_out = temp_data_out + shift_reg[279] * COEFF_279;
        temp_data_out = temp_data_out + shift_reg[280] * COEFF_280;
        temp_data_out = temp_data_out + shift_reg[281] * COEFF_281;
        temp_data_out = temp_data_out + shift_reg[282] * COEFF_282;
        temp_data_out = temp_data_out + shift_reg[283] * COEFF_283;
        temp_data_out = temp_data_out + shift_reg[284] * COEFF_284;
        temp_data_out = temp_data_out + shift_reg[285] * COEFF_285;
        temp_data_out = temp_data_out + shift_reg[286] * COEFF_286;
        temp_data_out = temp_data_out + shift_reg[287] * COEFF_287;
        temp_data_out = temp_data_out + shift_reg[288] * COEFF_288;
        temp_data_out = temp_data_out + shift_reg[289] * COEFF_289;
        temp_data_out = temp_data_out + shift_reg[290] * COEFF_290;
        temp_data_out = temp_data_out + shift_reg[291] * COEFF_291;
        temp_data_out = temp_data_out + shift_reg[292] * COEFF_292;
        temp_data_out = temp_data_out + shift_reg[293] * COEFF_293;
        temp_data_out = temp_data_out + shift_reg[294] * COEFF_294;
        temp_data_out = temp_data_out + shift_reg[295] * COEFF_295;
        temp_data_out = temp_data_out + shift_reg[296] * COEFF_296;
        temp_data_out = temp_data_out + shift_reg[297] * COEFF_297;
        temp_data_out = temp_data_out + shift_reg[298] * COEFF_298;
        temp_data_out = temp_data_out + shift_reg[299] * COEFF_299;
        temp_data_out = temp_data_out + shift_reg[300] * COEFF_300;
        temp_data_out = temp_data_out + shift_reg[301] * COEFF_301;
        temp_data_out = temp_data_out + shift_reg[302] * COEFF_302;
        temp_data_out = temp_data_out + shift_reg[303] * COEFF_303;
        temp_data_out = temp_data_out + shift_reg[304] * COEFF_304;
        temp_data_out = temp_data_out + shift_reg[305] * COEFF_305;
        temp_data_out = temp_data_out + shift_reg[306] * COEFF_306;
        temp_data_out = temp_data_out + shift_reg[307] * COEFF_307;
        temp_data_out = temp_data_out + shift_reg[308] * COEFF_308;
        temp_data_out = temp_data_out + shift_reg[309] * COEFF_309;
        temp_data_out = temp_data_out + shift_reg[310] * COEFF_310;
        temp_data_out = temp_data_out + shift_reg[311] * COEFF_311;
        temp_data_out = temp_data_out + shift_reg[312] * COEFF_312;
        temp_data_out = temp_data_out + shift_reg[313] * COEFF_313;
        temp_data_out = temp_data_out + shift_reg[314] * COEFF_314;
        temp_data_out = temp_data_out + shift_reg[315] * COEFF_315;
        temp_data_out = temp_data_out + shift_reg[316] * COEFF_316;
        temp_data_out = temp_data_out + shift_reg[317] * COEFF_317;
        temp_data_out = temp_data_out + shift_reg[318] * COEFF_318;
        temp_data_out = temp_data_out + shift_reg[319] * COEFF_319;
        temp_data_out = temp_data_out + shift_reg[320] * COEFF_320;
        temp_data_out = temp_data_out + shift_reg[321] * COEFF_321;
        temp_data_out = temp_data_out + shift_reg[322] * COEFF_322;
        temp_data_out = temp_data_out + shift_reg[323] * COEFF_323;
        temp_data_out = temp_data_out + shift_reg[324] * COEFF_324;
        temp_data_out = temp_data_out + shift_reg[325] * COEFF_325;
        temp_data_out = temp_data_out + shift_reg[326] * COEFF_326;
        temp_data_out = temp_data_out + shift_reg[327] * COEFF_327;
        temp_data_out = temp_data_out + shift_reg[328] * COEFF_328;
        temp_data_out = temp_data_out + shift_reg[329] * COEFF_329;
        temp_data_out = temp_data_out + shift_reg[330] * COEFF_330;
        temp_data_out = temp_data_out + shift_reg[331] * COEFF_331;
        temp_data_out = temp_data_out + shift_reg[332] * COEFF_332;
        temp_data_out = temp_data_out + shift_reg[333] * COEFF_333;
        temp_data_out = temp_data_out + shift_reg[334] * COEFF_334;
        temp_data_out = temp_data_out + shift_reg[335] * COEFF_335;

        // Update data_out at the end of accumulation using non-blocking assignment
        data_out <= temp_data_out;
    end
end

endmodule
